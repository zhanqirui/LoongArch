`define FS_TO_DS_WD 64
`define DS_TO_ES_WD 148
`define ES_TO_MS_WD 71
`define MS_TO_WS_WD 70

`define WS_TO_RF_WD 37

`define BR_TO_FS_WD 5
