`define FS_TO_DS_WD 64
`define DS_TO_ES_WD 148
`define ES_TO_MS_WD 71
`define MS_TO_WS_WD 70

`define WS_TO_RF_WD 38

`define BR_TO_FS_WD 33

`define DS_TO_CHE_WD 11

`define ES_TO_CHE_WD 6
`define MS_TO_CHE_WD 6
